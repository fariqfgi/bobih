module bobih

pub fn main() string {
   return $tmpl('../../../../../../flag')
}
